module char

fn test_chars_do_born() {
	one := init_character('one')
	two := init_character('two')
	println('one: $one, two: $two')
}